module keydetect(	input [7:0] keycode, keycode1, keycode2, keycode3, keycode4, keycode5, targetkeycode,
						output key_on
						);