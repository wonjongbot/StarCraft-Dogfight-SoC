module joystick	(	input logic clk,
							output logic [1:0] x, y,
							otuput logic [2:] button);